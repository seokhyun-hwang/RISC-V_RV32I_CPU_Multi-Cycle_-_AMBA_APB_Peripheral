`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:2**8-1];
    /*
    initial begin
       // $readmemh("code.mem", rom);
        
        //rom[x]=32'b   f7  _ rs2 _ rs1 _ f3_ rd  _ opcode;  // R-Type
        rom[0] = 32'b0000000_00001_00010_000_00100_0110011;  // add x4, x2, x1;
        rom[1] = 32'b0100000_00001_00010_000_00101_0110011;  // sub x5, x2, x1;
        rom[2] = 32'b0000000_00000_00011_111_00110_0110011;  // and x6, x3, x0;
        rom[3] = 32'b0000000_00000_00011_110_00111_0110011;  // or  x7, x3, x0;

        //rom[x]=32'b    imm     _ rs1 _ f3_ rd  _ opcode;  // I-Type
        rom[4] = 32'b000000000001_00001_000_01001_0010011;  // addi  x9, x1,  1;
        rom[5] = 32'b000000000100_00010_111_01010_0010011;  // andi x10, x2,  4;
        rom[6] = 32'b000000000011_00001_001_01011_0010011;  // slli x11, x1,  3;
        rom[7] = 32'b000000001001_00001_001_01100_0010011;  // slli x12, x1,  9;
        rom[8] = 32'b000000011110_00001_001_01101_0010011;  // slli x13, x1, 30;

        //rom[x]= 32'b imm7 _ rs2 _ rs1 _f3 _imm5 _ opcode;  // B-Type  
        rom[9] = 32'b0000000_00010_00010_000_01100_1100011;  // beq x2, x2, 12;

        //rom[x]= 32'b  imm  _ rs2 _ rs1 _f3 _ imm _ opcode;  // S-Type  
        rom[12] = 32'b0000000_01011_00000_000_00100_0100011;  // sb x11,  4(x0);
        rom[13] = 32'b0000000_01100_00000_001_01000_0100011;  // sh x12,  8(x0);
        rom[14] = 32'b0000000_01101_00000_010_01100_0100011;  // sw x13, 12(x0);

        //rom[x]= 32'b    imm     _ rs1 _f3 _ rd  _ opcode;  // L-Type  
        rom[15] = 32'b000000000100_00000_000_01110_0000011;  // lb x14,  4(x0);
        rom[16] = 32'b000000001000_00000_001_01111_0000011;  // lh x15,  8(x0);
        rom[17] = 32'b000000001100_00000_010_10000_0000011;  // lw x16, 12(x0);

        //rom[x]= 32'b        imm         _ rd  _ opcode;  // LU-Type  
        rom[18] = 32'b00010000000000000000_10001_0110111;  // lui x17, 0x10000000;

        //rom[x]= 32'b        imm         _ rd  _ opcode;  // AU-Type  
        rom[19] = 32'b00010000000000000000_10010_0010111;  // auipc x18, 0x10000000;

        //rom[x]= 32'b         imm        _ rd  _ opcode;  // J-Type  
        rom[20] = 32'b00000001000000000000_00011_1101111;  // jal x3, 16

        //rom[x]= 32'b    imm     _ rs1 _f3 _ rd  _ opcode;  // JL-Type  
        rom[24] = 32'b000000011100_00100_000_00100_1100111;  // jalr x4, 28(x4); 
    end*/

    // Testbench initial 블록에서 이 ROM을 초기화합니다.
    initial begin
        // nop (addi x0, x0, 0)
        logic [31:0] nop = 32'h00000013;

        // --- R-type (index 0-9) ---
        // (x1=1, x2=2, x3=3, x0=0 가정)
        rom[0] = 32'b0000000_00001_00010_000_00100_0110011;  // 0: add  x4, x2, x1   (x4 = 3)
        rom[1] = 32'b0100000_00001_00010_000_00101_0110011;  // 1: sub  x5, x2, x1   (x5 = 1)
        rom[2] = 32'b0000000_00000_00011_111_00110_0110011;  // 2: and  x6, x3, x0   (x6 = 0)
        rom[3] = 32'b0000000_00000_00011_110_00111_0110011;  // 3: or   x7, x3, x0   (x7 = 3)
        rom[4] = 32'b0000000_00010_00001_001_01000_0110011;  // 4: sll  x8, x1, x2   (x8 = 4)
        rom[5] = 32'b0000000_00010_00001_010_01001_0110011;  // 5: slt  x9, x1, x2   (x9 = 1)
        rom[6] = 32'b0000000_00010_00001_011_01010_0110011;  // 6: sltu x10, x1, x2  (x10 = 1)
        rom[7] = 32'b0000000_00010_00001_100_01011_0110011;  // 7: xor  x11, x1, x2  (x11 = 3)
        rom[8] = 32'b0000000_00010_00001_101_01100_0110011;  // 8: srl  x12, x1, x2  (x12 = 0)
        rom[9] = 32'b0100000_00010_00001_101_01101_0110011;  // 9: sra  x13, x1, x2  (x13 = 0)

        // --- I-type (Arithmetic) (index 10-18) ---
        rom[10] = 32'b000000000001_00001_000_01110_0010011;  // 10: addi  x14, x1, 1    (x14 = 2)
        rom[11] = 32'b000000000100_00010_111_01111_0010011;  // 11: andi  x15, x2, 4    (x15 = 0)
        rom[12] = 32'b000000000101_00001_010_10000_0010011;  // 12: slti  x16, x1, 5    (x16 = 1)
        rom[13] = 32'b000000000101_00001_011_10001_0010011;  // 13: sltiu x17, x1, 5    (x17 = 1)
        rom[14] = 32'b000000000101_00001_100_10010_0010011;  // 14: xori  x18, x1, 5    (x18 = 4)
        rom[15] = 32'b000000000101_00001_110_10011_0010011;  // 15: ori   x19, x1, 5    (x19 = 5)
        rom[16] = 32'b0000000_00011_00001_001_10100_0010011;  // 16: slli  x20, x1, 3    (x20 = 8)
        rom[17] = 32'b0000000_00010_00001_101_10101_0010011;  // 17: srli  x21, x1, 2    (x21 = 0)
        rom[18] = 32'b0100000_00010_00001_101_10110_0010011;  // 18: srai  x22, x1, 2    (x22 = 0)


        // --- [수정] S-type을 위한 값 준비 (x30 = 0xFFEEDDCC) (index 24-25) ---
        rom[24] = 32'hFFEEDF37;  // 24: lui x30, 0xFFEED (x30 = 0xFFEED000)
        rom[25] = 32'hDCCF0F13;  // 25: addi x30, x30, 0xDCC (x30 = 0xFFEEDDCC)
        // --- S-type [실행] (RAM 덮어쓰기) (index 26-28) ---
        // (x30 = 0xFFEEDDCC)
        rom[26] = 32'b0000000_11110_00000_000_10000_0100011; // 26: sb x30, 16(x0)  (MEM[16] = 0xCC)
        rom[27] = 32'b0000000_11110_00000_001_10100_0100011; // 27: sh x30, 20(x0)  (MEM[20:21] = 0xDDCC)
        rom[28] = 32'b0000000_11110_00000_010_11000_0100011; // 28: sw x30, 24(x0)  (MEM[24:27] = 0xFFEEDDCC)

        // --- L-type [Post-Check] (S-type 결과 읽기) (index 29-33) ---
        rom[29] = 32'b000000010000_00000_000_00100_0000011; // 29: lb  x4, 16(x0)   (x4 = 0xFFFFFFCC, 부호확장)
        rom[30] = 32'b000000010100_00000_001_00101_0000011; // 30: lh  x5, 20(x0)   (x5 = 0xFFFFDDCC, 부호확장)
        rom[31] = 32'b000000011000_00000_010_00110_0000011; // 31: lw  x6, 24(x0)   (x6 = 0xFFEEDDCC)
        rom[32] = 32'b000000010000_00000_100_00111_0000011; // 32: lbu x7, 16(x0)   (x7 = 0x000000CC, 제로확장)
        rom[33] = 32'b000000010100_00000_101_01000_0000011; // 33: lhu x8, 20(x0)   (x8 = 0x0000DDCC, 제로확장)

        // --- B-type (Branch) (index 27~) ---
        // 각 브랜치가 성공하면 3개의 nop를 건너뛰도록 offset = 16 (4 명령어)로 설정.

        // Test 1: beq (x1=1, x2=2, 1==2는 false -> No Branch)
        rom[30] = 32'b0000000_00010_00001_000_10000_1100011;  // 27: beq  x1, x2, 16 (No Branch)


        // Test 2: bne (x1=1, x2=2, 1!=2는 true -> Branch!)
        rom[31] = 32'b0000000_00010_00001_001_10000_1100011;  // 31: bne  x1, x2, 16 (Branch!)

        // PC가 35로 점프 (31*4 + 16 = 124 + 16 = 140. 140/4 = 35)

        // Test 3: blt (x1=1, x2=2, 1<2는 true -> Branch!)
        rom[35] = 32'b0000000_00010_00001_100_10000_1100011;  // 35: blt  x1, x2, 16 (Branch!)

        // PC가 39로 점프

        // Test 4: bge (x1=1, x2=2, 1>=2는 false -> No Branch)
        rom[39] = 32'b0000000_00010_00001_101_10000_1100011;  // 39: bge  x1, x2, 16 (No Branch)
        rom[40] = nop;  // 40: nop (Executed)
        rom[41] = nop;  // 41: nop (Executed)
        rom[42] = nop;  // 42: nop (Executed)

        // Test 5: bltu (x1=1, x2=2, 1<2는 true -> Branch!)
        rom[43] = 32'b0000000_00010_00001_110_10000_1100011;  // 43: bltu x1, x2, 16 (Branch!)

        // PC가 47로 점프

        // Test 6: bgeu (x1=1, x2=2, 1>=2는 false -> No Branch)
        rom[47] = 32'b0000000_00010_00001_111_10000_1100011;  // 47: bgeu x1, x2, 16 (No Branch)


        // --- U-type (index 51-52) ---
        rom[51] = 32'b00010000000000000000_11100_0110111; // 51: lui   x28, 0x10000 (x28 = 0x10000000)
        rom[52] = 32'b00010000000000000000_11101_0010111; // 52: auipc x29, 0x10000 (x29 = PC + 0x10000000)
                                                          // (PC = 52*4 = 208. x29 = 208 + 0x10000000)

        // --- J-type (JAL) (index 53) ---
        // 3개의 nop를 건너뛰도록 offset = 16 (4 명령어)로 설정.
        rom[53] = 32'b00000001000000000000_00011_1101111;  // 53: jal x3, 16 (x3=PC+4, PC=PC+16)
        rom[54] = nop;  // 54: nop (Skipped)
        rom[55] = nop;  // 55: nop (Skipped)
        rom[56] = nop;  // 56: nop (Skipped)
        // PC가 57로 점프 (53*4 + 16 = 212 + 16 = 228. 228/4 = 57)
        // x3 = 53*4 + 4 = 216

        // --- J-type (JALR) (index 57) ---
        // (x1=1) + 28 = 29. LSB가 0이 되어 28로 점프. (index 7)
        rom[57] = 32'b000000011100_00001_000_00100_1100111; // 57: jalr x4, 28(x1) (x4=PC+4, PC=x1+28)
        // PC가 7번 인덱스 (rom[7])로 점프.
        // x4 = 57*4 + 4 = 232

        // --- End ---
        // 나머지는 nop로 채움
        for (int i = 58; i < 64; i++) begin
            rom[i] = nop;
        end
    end


    assign data = rom[addr[31:2]];
endmodule
